/*
File: cordic_core.v
Modules: cordic_core
Heirarchy: cordic_core

Created : 28/2/2016

*/

/*
Module: cordic_core
*/

module cordic_core(
	clk,
	reset_n,


);
